library verilog;
use verilog.vl_types.all;
entity comp_8bits_tb is
end comp_8bits_tb;
